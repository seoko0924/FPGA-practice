`timescale 1ns / 1ps

module tb_alu;

    // 1. 입력 (값을 바꿔가며 테스트해야 하므로 reg)
    reg [3:0] a;
    reg [3:0] b;
    reg [1:0] op;

    // 2. 출력 (결과를 받아야 하므로 wire)
    wire [3:0] y;

    // 3. ALU 모듈 연결 (Unit Under Test)
    alu u1 (
        .a(a), 
        .b(b), 
        .op(op), 
        .y(y)
    );

    initial begin
        $display("=== ALU Simulation Start ===");
        // 시간, Op코드, 입력값(2진수/10진수), 결과값(2진수/10진수)을 실시간 감시
        $monitor("Time=%0t | Op=%b | A=%b(%d) B=%b(%d) | Result Y=%b(%d)", 
                 $time, op, a, a, b, b, y, y);

        // 초기값 설정
        a = 4'b1100; // 10진수 12
        b = 4'b1010; // 10진수 10
        op = 2'b00;
        #10;

        // ==========================================
        // Case 1: AND 연산 (Op = 00)
        // 1100 & 1010 = 1000 (8)
        // ==========================================
        op = 2'b00;
        #10;

        // ==========================================
        // Case 2: OR 연산 (Op = 01)
        // 1100 | 1010 = 1110 (14)
        // ==========================================
        op = 2'b01;
        #10;

        // ==========================================
        // Case 3: XOR 연산 (Op = 10)
        // 1100 ^ 1010 = 0110 (6)
        // ==========================================
        op = 2'b10;
        #10;

        // ==========================================
        // Case 4: 덧셈 연산 (Op = 11)
        // 12 + 10 = 22 (10110) 이지만 4비트라 잘림 -> 6 (0110)
        // ==========================================
        op = 2'b11;
        #10;

        // 덧셈 테스트 하나 더 (작은 수)
        // 3 + 2 = 5 (0101)
        a = 3; b = 2;
        #10;

        $display("=== Simulation Finish ===");
        $stop;
    end

endmodule