`timescale 1ns / 1ps



module tb_mux_2x1;

    reg d0;
    reg d1;
    reg sel;
    wire y;
    
    mux_2x1 u1(.d0(d0),.d1(d1),.sel(sel),.y(y));
    
    initial begin
        $display("=== Mux 2x1 Simulation Start ===");
        // 시간, 선택신호, 입력값들, 그리고 결과를 실시간으로 감시
        $monitor("Time=%0t | Sel=%b | d0=%b d1=%b | Output y=%b", 
                 $time, sel, d0, d1, y);

        // [초기화] 모든 입력 0으로 시작
        sel = 0; d0 = 0; d1 = 0;
        #10;

        // ==========================================
        // 시나리오 1: Sel = 0일 때 (d0가 통과해야 함)
        // ==========================================
        $display("-- Check Channel 0 (Sel=0) --");
        sel = 0;
        
        d0 = 1; d1 = 0; // d0만 1로 바꿈 -> y도 1이 되어야 함
        #10;
        
        d0 = 0; d1 = 1; // d1을 1로 바꿨지만 sel=0이라서 무시되어야 함 (y=0 유지)
        #10;

        // ==========================================
        // 시나리오 2: Sel = 1일 때 (d1이 통과해야 함)
        // ==========================================
        $display("-- Check Channel 1 (Sel=1) --");
        sel = 1;
        
        d0 = 1; d1 = 0; // d0가 1이지만 sel=1이라서 무시되어야 함 (y=0 유지)
        #10;
        
        d0 = 0; d1 = 1; // d1을 1로 바꿈 -> y도 1이 되어야 함
        #10;

        // ==========================================
        // 시나리오 3: 스위칭 테스트
        // ==========================================
        $display("-- Switching Test --");
        d0 = 1; d1 = 0; // d0는 1, d1은 0인 상태
        
        sel = 0; #10;   // y는 d0를 따라가니까 1
        sel = 1; #10;   // y는 d1을 따라가니까 0
        sel = 0; #10;   // 다시 1

        $display("=== Simulation Finish ===");
        $stop;
    end
endmodule
