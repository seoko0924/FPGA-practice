`timescale 1ns / 1ps


module d_flip_flop(
    input clk,
    input rst,
    input d,
    output reg q

    );
    always @(posedge clk or posedge  rst) begin
        if (rst) begin
            q <= 1'b0;
        end
        else q <= d;
    end
    
endmodule
